//立即数生成模块
// 修订历史 :
// --------------------------------------------------------------------
//   版本 | 作者  | 修改日期    | 所做改变
//   V1.0 | 233  | 2020.6.24   | 肖老师给的初始版本
//   v1.1 | 233  | 2020.6.26   | 增加S型立即数的生成  
//   v1.2 | 233  | 2020.6.26   | 增加J,U,B型立即数的生成  
// --------------------------------------------------------------------
module ImmeGen(
   input  logic [4:0] iImm_type,
   input  logic [31:0] iInstruction,
   output logic [31:0] oImmediate
);
   wire [31:0]  instr = iInstruction;     // 换一个短点的符号
   wire [31:0]  i_imm = { {20{instr[31]}}, instr[31:20] };  
   //符号位扩展的方法，高位补足符号位（也说明了RISC-V的立即数是有符号数）

   /***********   v1.1 | 233  | 2020.6.26   | 增加S型立即数的生成  ***********/
   wire [31:0]  s_imm = { {20{instr[31]}} , instr[31:25] , instr[11:7] };
   /*************************************************************************/


   /**********v1.2 | 233  | 2020.6.26   | 增加J,U,B型立即数的生成  **********/
   logic tool_zero;              //工具数0
   assign tool_zero = 1'b0;
   wire [31:0]  b_imm = { {19{instr[31]}},instr[31],instr[7],
                           instr[30:25],instr[11:8],tool_zero };

   wire [31:0]  u_imm = { instr[31:12] , { 12{tool_zero} } };

   wire [31:0]  j_imm = { {11{tool_zero}} , instr[31] , instr[19:12] , instr[20] , 
                           instr[30:21] , tool_zero };
   /*************************************************************************/


   // 使用与或门的方法构成多路数据选择器
   wire iJ_type, iU_type, iB_type, iS_type, iI_type;  //立即数类型信号
   assign {iJ_type, iU_type, iB_type, iS_type, iI_type} = iImm_type;
                                                      //传递立即数类型信号，确定立即数类型
   assign  oImmediate = ({32{iI_type}} & i_imm)
   
   /******************   v1.1 | 233  | 2020.6.26   | 增加S型立即数的生成  ******************/   
                        | ({32{iS_type}} & s_imm)
   /**************************************************************************************/
   
   /**********v1.2 | 233  | 2020.6.26   | 增加J,U,B型立即数的生成  **********/
                        | ({32{iB_type}} & b_imm)
                        | ({32{iU_type}} & u_imm)
                        | ({32{iJ_type}} & j_imm)
      ;
   /*************************************************************************/
endmodule
